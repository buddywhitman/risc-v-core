module inst_mem(
	input clk,
	input [31:0] addr,
	output [31:0] read_data
);
	reg [31:0] mem [0 : 31];
	assign read_data = mem[addr];
	
	always @(posedge clk)
	begin
		mem[0] = {32{1'b0}};
		mem[1] = 32'b000000000011_00000_000_00101_0010011;
		mem[2] = 32'b000000000101_00000_000_00110_0010011;
		mem[3] = 32'b000000000110_00101_000_00111_0110011;
		mem[4] = 32'b00000000011100000_010_00011_0100011;
		mem[5] = 32'b11111110101001000010101000100011;
		mem[6] = 32'b11111111010001000010010100000011;
		mem[7] = 32'b00000000101001010000010100110011;
		mem[8] = 32'b00000000100000010010010000000011;
		mem[9] = 32'b00000000110000010010000010000011;
		mem[10] = 32'b00000001000000010000000100010011;
		mem[11] = 32'b00000000000000001000000001100111;
		
	
	end
endmodule
